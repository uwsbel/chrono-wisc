!!!! CIURCUIT !!!!
RaC n5 n1 {parRaC}
LaC n4 n5 {parLaC} ic{icLaC}
VbackemfCVAR n4 n3 PWL(0 0 1e-9 0)
Vprobe1 n2 n3 0
VgenVAR n6 0 PWL(0 0 1e-9 0)
S1 n12 n6 n10 0 SW1
VSW1VAR n10 0 PWL(0 0 1e-9 0)
X1 n1 n8 n7 irf520
D1 n1 n2 DI_1N4007
C1 n2 n11 12e-6
R8 n11 n1 25
R1 n7 0 2
R3 n12 n2 15
VgenPWMVAR n8 0 PWL(0 0 1e-9 0)
R2 n8 0 10e3
VMos1 n9 0 25
.param parVgenVAR=0.0
.param parVbackemfCVAR=0.0
.param parLaC=45.0e-6
.param parRaC=25.1
.param parVSW1VAR=0.0
.param parVgenPWMVAR=0.0
.param icLaC=0.000000e+00
.ic 
**********MODELS**********
*****MODEL1*****
.model SW1 SW(Ron=0.1 Roff=1Meg Vt=.5 Vh=0)
*****MODEL2*****
.MODEL DI_1N4007 D  ( IS=76.9p RS=42.0m BV=1.00k IBV=5.00u
+ CJO=26.5p  M=0.333 N=1.45 TT=4.32u )
*****MODEL3*****
.SUBCKT irf520 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.61397 LAMBDA=0.00572642 KP=3.9143
+CGSO=3.28344e-06 CGDO=1.0112e-11
RS 8 3 0.171045
D1 3 1 MD
.MODEL MD D IS=7.10668e-11 RS=0.0302634 N=1.21428 BV=100
+IBV=0.00025 EG=1 XTI=2.99378 TT=2.27818e-09
+CJO=5.01988e-10 VJ=0.565258 M=0.378444 FC=0.5
RDS 3 1 4e+06
RD 9 1 0.01473
RG 2 7 1.34402
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=4.14565e-10 VJ=0.5 M=0.640575 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=1e-10 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 6.23795e-10
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.4
.ENDS